module Battleship;


endmodule
