module contar_unos_operador(input [4:0] numero, output [3:0] cantidad_unos);
    logic[4:0] unos;

	assign cantidad_unos = unos;
	
	always @(numero)
	begin
		case(numero)
		// 0000 -> 0
		5'b00000:unos = 4'b0000;
		
		// 0001 -> 1 
		5'b00001: unos = 4'b0001;
		
		// 0010 -> 2
		5'b00010: unos = 4'b0001;
		
		// 0011 -> 3 
		5'b00011: unos = 4'b0010;
		
		// 0100 -> 4
		5'b00100: unos = 4'b0001;
		
		// 0101 -> 5 
		5'b00101: unos = 4'b0010;
		
		// 0110 -> 6
		5'b00110: unos = 4'b0010;
		
		// 0111 -> 7 
		5'b00111: unos = 4'b0011;
	
		// 1000 -> 8
		5'b01000: unos = 4'b0001;
		
		// 1001 -> 9 
		5'b01001: unos = 4'b0010;
		
		// 1010 -> 10 
		5'b01010: unos = 4'b0010;
		
		// 01011 -> 11 
		5'b01011: unos = 4'b0011;
		
		// 01100 -> 12
		5'b01100: unos = 4'b0010;
		
		// 01101 -> 13 
		5'b01101: unos = 4'b0011;
		
		// 01110 -> 14 
		5'b01110: unos = 4'b0011;
		
		// 01111 -> 15 
		5'b01111: unos = 4'b0100;
		
		// 10000 -> 16
		5'b10000:unos = 4'b0001;
		
		// 0001 -> 17 
		5'b10001: unos = 4'b0010;
		
		// 10010 -> 18
		5'b10010: unos = 4'b0010;
		
		// 10011 -> 19 
		5'b10011: unos = 4'b0011;
		
		// 10100 -> 20
		5'b10100: unos = 4'b0010;
		
		// 10101 -> 21 
		5'b10101: unos = 4'b0011;
		
		// 10110 -> 22
		5'b10110: unos = 4'b0011;
		
		// 10111 -> 23 
		5'b10111: unos = 4'b0100;
	
		// 11000 -> 24
		5'b11000: unos = 4'b0010;
		
		// 11001 -> 25 
		5'b11001: unos = 4'b0011;
		
		// 11010 -> 26 
		5'b11010: unos = 4'b0011;
		
		// 11011 -> 27 
		5'b11011: unos = 4'b0100;
		
		// 11100 -> 28
		5'b11100: unos = 4'b0011;
		
		// 11101 -> 29 
		5'b11101: unos = 4'b0100;
		
		// 11110 -> 30 
		5'b11110: unos = 4'b0100;
		
		// 11111 -> 31 
		5'b11111: unos = 4'b0101;
		
		endcase
	end
endmodule
