module divider_8bit(
  input logic [7:0] dividend,
  input logic [7:0] divisor,
  output logic [7:0] quotient,
  output logic overflow,
  output logic zero
  
);

  

endmodule